{"File":{"Name":"03-02T03:35:17_52a8_W037","Program":"BEATmonitor/survey","Version":"v0.01","Firmware":"2v25","Serial":"963a869d-d057e561","MAC":"d8:8a:52:0a:52:a8","PhysicalID":"W037"}}
null
{"timeStamp":1740880951290.96215820312,"question":"FAMILIAR","input":"slider","range":[0,6],"response":"NA"}
{"timeStamp":1740886517629.34106445312,"question":"LIKE","input":"slider","range":[0,6],"response":"NA"}