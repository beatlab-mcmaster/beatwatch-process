{"File":{"Name":"03-02T01:53:40_f937_W025","Program":"BEATmonitor/survey","Version":"v0.01","Firmware":"2v25","Serial":"c915e4b8-57cc43fc","MAC":"e4:db:81:62:f9:37","PhysicalID":"W025"}}
{"Record":{"State":"START_RECORD","DateTime":"Sat Mar 1 2025 20:53:40 GMT-0500","UNIXTimeStamp":"2025-03-02T01:53:40.996Z","BatteryLife":76,"FreeStorage":4319692,"SamplesWritten":0}}
{"timeStamp":1740880946410.61889648437,"question":"FAMILIAR","input":"slider","range":[0,6],"response":0}
{"timeStamp":1740880950862.76733398437,"question":"LIKE","input":"slider","range":[0,6],"response":2}
{"timeStamp":1740881047324.07104492187,"question":"FAMILIAR","input":"slider","range":[0,6],"response":6}
{"timeStamp":1740881057596.25732421875,"question":"LIKE","input":"slider","range":[0,6],"response":6}
{"timeStamp":1740881264887.24243164062,"question":"FAMILIAR","input":"slider","range":[0,6],"response":"NA"}
{"timeStamp":1740881269892.85766601562,"question":"LIKE","input":"slider","range":[0,6],"response":6}
{"timeStamp":1740882224402.5927734375,"question":"FAMILIAR","input":"slider","range":[0,6],"response":0}
{"timeStamp":1740882227532.7197265625,"question":"LIKE","input":"slider","range":[0,6],"response":3}
{"timeStamp":1740882482571.59912109375,"question":"FAMILIAR","input":"slider","range":[0,6],"response":6}
{"timeStamp":1740882491226.65893554687,"question":"LIKE","input":"slider","range":[0,6],"response":6}
{"timeStamp":1740882640741.73461914062,"question":"FAMILIAR","input":"slider","range":[0,6],"response":6}
{"timeStamp":1740882647357.64038085937,"question":"LIKE","input":"slider","range":[0,6],"response":6}
{"timeStamp":1740883758186.162109375,"question":"FAMILIAR","input":"slider","range":[0,6],"response":6}
{"timeStamp":1740883761773.35083007812,"question":"LIKE","input":"slider","range":[0,6],"response":6}
{"timeStamp":1740883794301.48803710937,"question":"FAMILIAR","input":"slider","range":[0,6],"response":6}
{"timeStamp":1740883799299.16870117187,"question":"LIKE","input":"slider","range":[0,6],"response":3}
{"Record":{"State":"STOP_RECORD","DateTime":"Sat Mar 1 2025 21:57:47 GMT-0500","UNIXTimeStamp":"2025-03-02T02:57:47.572Z","BatteryLife":77,"FreeStorage":1944012,"SamplesWritten":90985}}